*** Esempio scemo come la merda ***

vi n1 0 dc 1V ac 0V
R1 n3 n1 2.4k
C1 n3 0 2nF
.dc vi 0 100 0.01
.end
