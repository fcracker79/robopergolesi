*** Test NPN Inverter ***
*** plot v(pe)
.MODEL Q_NPN NPN(IS=800.0E-18 BF=2.000E3)
vi pin 0 dc 1V ac 0V
Q1 pe pb 0 Q_NPN
Re p2 pe 1k
Rb pin pb 20k
vl p2 0 dc 4.8V ac 0V
.dc vi -1.5 1.5 0.01
.end
